// inputs:
//
// outputs:
//
module ethernet_controller ;

endmodule // ethernet_controller
