library verilog;
use verilog.vl_types.all;
entity ProtocolInfo is
end ProtocolInfo;
