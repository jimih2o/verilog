library verilog;
use verilog.vl_types.all;
entity dm9000a_sv_unit is
end dm9000a_sv_unit;
